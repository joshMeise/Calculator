library IEEE;
use IEEE.std_logic_1164.all;

package myPackage is
  type opType is (sum, mult, sub);
end myPackage;
